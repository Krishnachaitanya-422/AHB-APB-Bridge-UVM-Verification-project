//abh agent