// virtual sequence