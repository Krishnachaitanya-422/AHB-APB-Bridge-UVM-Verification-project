//amba_vtest_lib