//ahb driver