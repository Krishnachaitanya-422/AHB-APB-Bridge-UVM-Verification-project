// top module

module top;
    
    import amba_test_pkg::*;
    import uvm_pkg::*;

    bit clk;

    
endmodule