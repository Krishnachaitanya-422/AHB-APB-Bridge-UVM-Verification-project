// ahb to apb env file