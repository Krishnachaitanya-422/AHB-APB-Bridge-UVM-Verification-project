//env config file