// top module