//test package file