//ahb monitor