//abh transaction