//abh transaction

class abh_trxn extends uvm_sequence_item;

	`uvm_object_utils(ahb_trxn)
	
	//Inputs and outputs:
	
	
	
	//Constraints
	
	
	
	extern function void do_print(uvm_printer printer);
endclass

/////----Constructor----/////

function void abh_trxn::do_print(uvm_printer printer);
		super.do_print(printer);
		
		
		//print statements
		
endfunction