//apb transaction

class apb_trxn extends uvm_sequence_item;
	
	`uvm_object_utils(apb_trxn)
	
	//I/p and O/P's
	
	
	
	//constraints


	extern function void do_print(uvm_printer);
	
	
endclass

function void apb_trxn::do_print(uvm_printer printer);
		super.do_print();
		
		//print statements
		
endfunction

