//ahb sequencer