//abh seqs