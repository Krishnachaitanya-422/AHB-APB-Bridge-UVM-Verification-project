//ahb agent top