//ahb agent config