// virtual sequencer